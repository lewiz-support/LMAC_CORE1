library verilog;
use verilog.vl_types.all;
entity tcore_fmac_core is
    generic(
        FMAC_ID         : integer := 10;
        RX_FIFO_DEPTH   : integer := 4096;
        RX_FIFO_ADDR_WIDTH: integer := 12;
        RX_DRAM_DEPTH   : integer := 3072;
        RX_DRAM_ADDR_WIDTH: integer := 12;
        OVERSIZE_MARK   : integer := 9022
    );
    port(
        usr_clk         : in     vl_logic;
        xaui_clk        : in     vl_logic;
        \usr_rst_\      : in     vl_logic;
        fmac_speed      : in     vl_logic_vector(1 downto 0);
        TCORE_MODE      : in     vl_logic;
        tx_xo_en        : in     vl_logic;
        rx_xo_en        : in     vl_logic;
        bcast_en        : in     vl_logic;
        prom_mode       : in     vl_logic;
        mac_addr0       : in     vl_logic_vector(47 downto 0);
        rx_size         : in     vl_logic_vector(11 downto 0);
        rx_check_crc    : in     vl_logic;
        txfifo_din      : in     vl_logic_vector(63 downto 0);
        txfifo_wr_en    : in     vl_logic;
        txfifo_full     : out    vl_logic;
        txfifo_usedw    : out    vl_logic_vector(12 downto 0);
        mac_pause_value : in     vl_logic_vector(31 downto 0);
        tx_b2b_dly      : in     vl_logic_vector(1 downto 0);
        rxfifo_rd_cycle : in     vl_logic;
        rxfifo_rd_en    : in     vl_logic;
        rxfifo_dout     : out    vl_logic_vector(63 downto 0);
        rxfifo_ctrl_dout: out    vl_logic_vector(7 downto 0);
        rxfifo_empty    : out    vl_logic;
        rxfifo_full_dbg : out    vl_logic;
        rxfifo_usedw_dbg: out    vl_logic_vector;
        drx_pkt_data    : out    vl_logic_vector(63 downto 0);
        drx_pkt_start   : out    vl_logic;
        drx_pkt_end     : out    vl_logic;
        drx_pkt_we      : out    vl_logic;
        drx_pkt_beat_bcnt: out    vl_logic_vector(2 downto 0);
        drx_pkt_be      : out    vl_logic_vector(7 downto 0);
        drx_crc32       : out    vl_logic_vector(31 downto 0);
        drx_crc_vld     : out    vl_logic;
        drx_crc_err     : out    vl_logic;
        drx_crc_err_dly1: out    vl_logic;
        cs_fifo_rd_en   : in     vl_logic;
        ipcs_fifo_dout  : out    vl_logic_vector(63 downto 0);
        cs_fifo_empty   : out    vl_logic;
        xgmii_rxc       : in     vl_logic_vector(7 downto 0);
        xgmii_rxd       : in     vl_logic_vector(63 downto 0);
        xgmii_rxp       : in     vl_logic_vector(7 downto 0);
        br_sof4         : in     vl_logic;
        fmac_ctrl1_dly  : in     vl_logic_vector(31 downto 0);
        fmac_rxd_en     : in     vl_logic;
        gmii_txd        : out    vl_logic_vector(7 downto 0);
        gmii_txc        : out    vl_logic;
        gmii_tx_en      : out    vl_logic;
        gmii_tx_vld     : out    vl_logic;
        linkup_1g       : in     vl_logic;
        gige_clk        : in     vl_logic;
        FMAC_TX_PKT_CNT : out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT_LO: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT_HI: out    vl_logic_vector(31 downto 0);
        FMAC_TX_BYTE_CNT: out    vl_logic_vector(31 downto 0);
        FMAC_RX_BYTE_CNT_LO: out    vl_logic_vector(31 downto 0);
        FMAC_RX_BYTE_CNT_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_UNDERSIZE_PKT_CNT: out    vl_logic_vector(31 downto 0);
        FMAC_RX_CRC_ERR_CNT: out    vl_logic_vector(31 downto 0);
        FMAC_DCNT_OVERRUN: out    vl_logic_vector(31 downto 0);
        FMAC_DCNT_LINK_ERR: out    vl_logic_vector(31 downto 0);
        FMAC_PKT_CNT_OVERSIZE: out    vl_logic_vector(31 downto 0);
        FIFO_OV_IPEND   : out    vl_logic;
        FMAC_PKT_CNT_JABBER: out    vl_logic_vector(31 downto 0);
        FMAC_PKT_CNT_FRAGMENT: out    vl_logic_vector(31 downto 0);
        STAT_GROUP_LO_DOUT: out    vl_logic_vector(31 downto 0);
        STAT_GROUP_HI_DOUT: out    vl_logic_vector(31 downto 0);
        STAT_GROUP_addr : in     vl_logic_vector(9 downto 0);
        STAT_GROUP_sel  : in     vl_logic;
        fmac_rx_clr_en  : in     vl_logic;
        fmac_tx_clr_en  : in     vl_logic;
        FMAC_RX_PKT_CNT64_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT64_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT127_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT127_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT255_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT255_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT511_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT511_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT1023_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT1023_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT1518_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT1518_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT2047_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT2047_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT4095_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT4095_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT8191_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT8191_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT9018_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT9018_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT9022_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT9022_HI: out    vl_logic_vector(31 downto 0);
        FMAC_RX_PKT_CNT9199P_LO: out    vl_logic_vector(32 downto 0);
        FMAC_RX_PKT_CNT9199P_HI: out    vl_logic_vector(31 downto 0)
    );
end tcore_fmac_core;
